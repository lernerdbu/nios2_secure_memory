// nios2_secure_memory.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module nios2_secure_memory (
		input  wire       clk_clk,                            //                         clk.clk
		output wire [7:0] led_pio_external_connection_export, // led_pio_external_connection.export
		input  wire       reset_reset_n                       //                       reset.reset_n
	);

	wire  [31:0] cpu_custom_instruction_master_result;                                  // cpu_custom_instruction_master_translator:ci_slave_result -> cpu:E_ci_combo_result
	wire         cpu_custom_instruction_master_readra;                                  // cpu:E_ci_combo_readra -> cpu_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] cpu_custom_instruction_master_a;                                       // cpu:E_ci_combo_a -> cpu_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] cpu_custom_instruction_master_b;                                       // cpu:E_ci_combo_b -> cpu_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] cpu_custom_instruction_master_c;                                       // cpu:E_ci_combo_c -> cpu_custom_instruction_master_translator:ci_slave_c
	wire         cpu_custom_instruction_master_readrb;                                  // cpu:E_ci_combo_readrb -> cpu_custom_instruction_master_translator:ci_slave_readrb
	wire         cpu_custom_instruction_master_estatus;                                 // cpu:E_ci_combo_estatus -> cpu_custom_instruction_master_translator:ci_slave_estatus
	wire  [31:0] cpu_custom_instruction_master_ipending;                                // cpu:E_ci_combo_ipending -> cpu_custom_instruction_master_translator:ci_slave_ipending
	wire  [31:0] cpu_custom_instruction_master_datab;                                   // cpu:E_ci_combo_datab -> cpu_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] cpu_custom_instruction_master_dataa;                                   // cpu:E_ci_combo_dataa -> cpu_custom_instruction_master_translator:ci_slave_dataa
	wire         cpu_custom_instruction_master_writerc;                                 // cpu:E_ci_combo_writerc -> cpu_custom_instruction_master_translator:ci_slave_writerc
	wire   [7:0] cpu_custom_instruction_master_n;                                       // cpu:E_ci_combo_n -> cpu_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] cpu_custom_instruction_master_translator_comb_ci_master_result;        // cpu_custom_instruction_master_comb_xconnect:ci_slave_result -> cpu_custom_instruction_master_translator:comb_ci_master_result
	wire         cpu_custom_instruction_master_translator_comb_ci_master_readra;        // cpu_custom_instruction_master_translator:comb_ci_master_readra -> cpu_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] cpu_custom_instruction_master_translator_comb_ci_master_a;             // cpu_custom_instruction_master_translator:comb_ci_master_a -> cpu_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] cpu_custom_instruction_master_translator_comb_ci_master_b;             // cpu_custom_instruction_master_translator:comb_ci_master_b -> cpu_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         cpu_custom_instruction_master_translator_comb_ci_master_readrb;        // cpu_custom_instruction_master_translator:comb_ci_master_readrb -> cpu_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] cpu_custom_instruction_master_translator_comb_ci_master_c;             // cpu_custom_instruction_master_translator:comb_ci_master_c -> cpu_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         cpu_custom_instruction_master_translator_comb_ci_master_estatus;       // cpu_custom_instruction_master_translator:comb_ci_master_estatus -> cpu_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] cpu_custom_instruction_master_translator_comb_ci_master_ipending;      // cpu_custom_instruction_master_translator:comb_ci_master_ipending -> cpu_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] cpu_custom_instruction_master_translator_comb_ci_master_datab;         // cpu_custom_instruction_master_translator:comb_ci_master_datab -> cpu_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] cpu_custom_instruction_master_translator_comb_ci_master_dataa;         // cpu_custom_instruction_master_translator:comb_ci_master_dataa -> cpu_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         cpu_custom_instruction_master_translator_comb_ci_master_writerc;       // cpu_custom_instruction_master_translator:comb_ci_master_writerc -> cpu_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] cpu_custom_instruction_master_translator_comb_ci_master_n;             // cpu_custom_instruction_master_translator:comb_ci_master_n -> cpu_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_result;         // cpu_custom_instruction_master_comb_slave_translator0:ci_slave_result -> cpu_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master0_readra;         // cpu_custom_instruction_master_comb_xconnect:ci_master0_readra -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_a;              // cpu_custom_instruction_master_comb_xconnect:ci_master0_a -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_b;              // cpu_custom_instruction_master_comb_xconnect:ci_master0_b -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb;         // cpu_custom_instruction_master_comb_xconnect:ci_master0_readrb -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_c;              // cpu_custom_instruction_master_comb_xconnect:ci_master0_c -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus;        // cpu_custom_instruction_master_comb_xconnect:ci_master0_estatus -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending;       // cpu_custom_instruction_master_comb_xconnect:ci_master0_ipending -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_datab;          // cpu_custom_instruction_master_comb_xconnect:ci_master0_datab -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa;          // cpu_custom_instruction_master_comb_xconnect:ci_master0_dataa -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc;        // cpu_custom_instruction_master_comb_xconnect:ci_master0_writerc -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_n;              // cpu_custom_instruction_master_comb_xconnect:ci_master0_n -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] cpu_custom_instruction_master_comb_slave_translator0_ci_master_result; // custom_secure_mem_instructions:result -> cpu_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab;  // cpu_custom_instruction_master_comb_slave_translator0:ci_master_datab -> custom_secure_mem_instructions:datab
	wire  [31:0] cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa;  // cpu_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> custom_secure_mem_instructions:dataa
	wire   [2:0] cpu_custom_instruction_master_comb_slave_translator0_ci_master_n;      // cpu_custom_instruction_master_comb_slave_translator0:ci_master_n -> custom_secure_mem_instructions:n
	wire         custom_secure_mem_instructions_avalon_master_chipselect;               // custom_secure_mem_instructions:chipselect -> mm_interconnect_0:custom_secure_mem_instructions_avalon_master_chipselect
	wire  [31:0] custom_secure_mem_instructions_avalon_master_readdata;                 // mm_interconnect_0:custom_secure_mem_instructions_avalon_master_readdata -> custom_secure_mem_instructions:readdata
	wire         custom_secure_mem_instructions_avalon_master_waitrequest;              // mm_interconnect_0:custom_secure_mem_instructions_avalon_master_waitrequest -> custom_secure_mem_instructions:waitrequest
	wire  [31:0] custom_secure_mem_instructions_avalon_master_address;                  // custom_secure_mem_instructions:address -> mm_interconnect_0:custom_secure_mem_instructions_avalon_master_address
	wire   [3:0] custom_secure_mem_instructions_avalon_master_byteenable;               // custom_secure_mem_instructions:byteenable -> mm_interconnect_0:custom_secure_mem_instructions_avalon_master_byteenable
	wire  [31:0] custom_secure_mem_instructions_avalon_master_writedata;                // custom_secure_mem_instructions:writedata -> mm_interconnect_0:custom_secure_mem_instructions_avalon_master_writedata
	wire         custom_secure_mem_instructions_avalon_master_write;                    // custom_secure_mem_instructions:write -> mm_interconnect_0:custom_secure_mem_instructions_avalon_master_write
	wire         mm_interconnect_0_onchip_mem_s2_chipselect;                            // mm_interconnect_0:onchip_mem_s2_chipselect -> onchip_mem:chipselect2
	wire  [31:0] mm_interconnect_0_onchip_mem_s2_readdata;                              // onchip_mem:readdata2 -> mm_interconnect_0:onchip_mem_s2_readdata
	wire  [12:0] mm_interconnect_0_onchip_mem_s2_address;                               // mm_interconnect_0:onchip_mem_s2_address -> onchip_mem:address2
	wire   [3:0] mm_interconnect_0_onchip_mem_s2_byteenable;                            // mm_interconnect_0:onchip_mem_s2_byteenable -> onchip_mem:byteenable2
	wire         mm_interconnect_0_onchip_mem_s2_write;                                 // mm_interconnect_0:onchip_mem_s2_write -> onchip_mem:write2
	wire  [31:0] mm_interconnect_0_onchip_mem_s2_writedata;                             // mm_interconnect_0:onchip_mem_s2_writedata -> onchip_mem:writedata2
	wire         mm_interconnect_0_onchip_mem_s2_clken;                                 // mm_interconnect_0:onchip_mem_s2_clken -> onchip_mem:clken2
	wire  [31:0] cpu_data_master_readdata;                                              // mm_interconnect_1:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                           // mm_interconnect_1:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                           // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:cpu_data_master_debugaccess
	wire  [16:0] cpu_data_master_address;                                               // cpu:d_address -> mm_interconnect_1:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                            // cpu:d_byteenable -> mm_interconnect_1:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                  // cpu:d_read -> mm_interconnect_1:cpu_data_master_read
	wire         cpu_data_master_write;                                                 // cpu:d_write -> mm_interconnect_1:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                             // cpu:d_writedata -> mm_interconnect_1:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                       // mm_interconnect_1:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                    // mm_interconnect_1:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [16:0] cpu_instruction_master_address;                                        // cpu:i_address -> mm_interconnect_1:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                           // cpu:i_read -> mm_interconnect_1:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                                  // mm_interconnect_1:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;              // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;                // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;             // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;                 // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;                    // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;                   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;               // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                        // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                         // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_cpu_debug_mem_slave_readdata;                        // cpu:debug_mem_slave_readdata -> mm_interconnect_1:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_1_cpu_debug_mem_slave_waitrequest;                     // cpu:debug_mem_slave_waitrequest -> mm_interconnect_1:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_1_cpu_debug_mem_slave_debugaccess;                     // mm_interconnect_1:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_1_cpu_debug_mem_slave_address;                         // mm_interconnect_1:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_1_cpu_debug_mem_slave_read;                            // mm_interconnect_1:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_1_cpu_debug_mem_slave_byteenable;                      // mm_interconnect_1:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_1_cpu_debug_mem_slave_write;                           // mm_interconnect_1:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_1_cpu_debug_mem_slave_writedata;                       // mm_interconnect_1:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_1_sys_clk_timer_s1_chipselect;                         // mm_interconnect_1:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_readdata;                           // sys_clk_timer:readdata -> mm_interconnect_1:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_1_sys_clk_timer_s1_address;                            // mm_interconnect_1:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_1_sys_clk_timer_s1_write;                              // mm_interconnect_1:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_writedata;                          // mm_interconnect_1:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_1_led_pio_s1_chipselect;                               // mm_interconnect_1:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_1_led_pio_s1_readdata;                                 // led_pio:readdata -> mm_interconnect_1:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_led_pio_s1_address;                                  // mm_interconnect_1:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_1_led_pio_s1_write;                                    // mm_interconnect_1:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_1_led_pio_s1_writedata;                                // mm_interconnect_1:led_pio_s1_writedata -> led_pio:writedata
	wire         mm_interconnect_1_onchip_mem_s1_chipselect;                            // mm_interconnect_1:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	wire  [31:0] mm_interconnect_1_onchip_mem_s1_readdata;                              // onchip_mem:readdata -> mm_interconnect_1:onchip_mem_s1_readdata
	wire  [12:0] mm_interconnect_1_onchip_mem_s1_address;                               // mm_interconnect_1:onchip_mem_s1_address -> onchip_mem:address
	wire   [3:0] mm_interconnect_1_onchip_mem_s1_byteenable;                            // mm_interconnect_1:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	wire         mm_interconnect_1_onchip_mem_s1_write;                                 // mm_interconnect_1:onchip_mem_s1_write -> onchip_mem:write
	wire  [31:0] mm_interconnect_1_onchip_mem_s1_writedata;                             // mm_interconnect_1:onchip_mem_s1_writedata -> onchip_mem:writedata
	wire         mm_interconnect_1_onchip_mem_s1_clken;                                 // mm_interconnect_1:onchip_mem_s1_clken -> onchip_mem:clken
	wire         irq_mapper_receiver0_irq;                                              // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                              // sys_clk_timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                                           // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                                        // rst_controller:reset_out -> [cpu:reset_n, irq_mapper:reset, mm_interconnect_1:cpu_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_reset_out_reset_req;                                    // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                                         // cpu:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                                    // rst_controller_001:reset_out -> [custom_secure_mem_instructions:reset, jtag_uart:rst_n, led_pio:reset_n, mm_interconnect_0:custom_secure_mem_instructions_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_reset_reset_bridge_in_reset_reset, onchip_mem:reset, onchip_mem:reset2, rst_translator_001:in_reset, sys_clk_timer:reset_n, sysid:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                                // rst_controller_001:reset_req -> [onchip_mem:reset_req, onchip_mem:reset_req2, rst_translator_001:reset_req_in]

	nios2_secure_memory_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_cpu_debug_mem_slave_writedata),   //                          .writedata
		.E_ci_combo_result                   (cpu_custom_instruction_master_result),              // custom_instruction_master.result
		.E_ci_combo_a                        (cpu_custom_instruction_master_a),                   //                          .a
		.E_ci_combo_b                        (cpu_custom_instruction_master_b),                   //                          .b
		.E_ci_combo_c                        (cpu_custom_instruction_master_c),                   //                          .c
		.E_ci_combo_dataa                    (cpu_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_combo_datab                    (cpu_custom_instruction_master_datab),               //                          .datab
		.E_ci_combo_estatus                  (cpu_custom_instruction_master_estatus),             //                          .estatus
		.E_ci_combo_ipending                 (cpu_custom_instruction_master_ipending),            //                          .ipending
		.E_ci_combo_n                        (cpu_custom_instruction_master_n),                   //                          .n
		.E_ci_combo_readra                   (cpu_custom_instruction_master_readra),              //                          .readra
		.E_ci_combo_readrb                   (cpu_custom_instruction_master_readrb),              //                          .readrb
		.E_ci_combo_writerc                  (cpu_custom_instruction_master_writerc)              //                          .writerc
	);

	secure_memory_top #(
		.xor_key (34'b0010010101110110100100111010101011)
	) custom_secure_mem_instructions (
		.dataa       (cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.datab       (cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //                              .datab
		.n           (cpu_custom_instruction_master_comb_slave_translator0_ci_master_n),      //                              .n
		.clk_en      (),                                                                      //                              .clk_en
		.start       (),                                                                      //                              .start
		.done        (),                                                                      //                              .done
		.result      (cpu_custom_instruction_master_comb_slave_translator0_ci_master_result), //                              .result
		.readdata    (custom_secure_mem_instructions_avalon_master_readdata),                 //                 avalon_master.readdata
		.address     (custom_secure_mem_instructions_avalon_master_address),                  //                              .address
		.writedata   (custom_secure_mem_instructions_avalon_master_writedata),                //                              .writedata
		.byteenable  (custom_secure_mem_instructions_avalon_master_byteenable),               //                              .byteenable
		.chipselect  (custom_secure_mem_instructions_avalon_master_chipselect),               //                              .chipselect
		.write       (custom_secure_mem_instructions_avalon_master_write),                    //                              .write
		.waitrequest (custom_secure_mem_instructions_avalon_master_waitrequest),              //                              .waitrequest
		.clk         (clk_clk),                                                               //                    clock_sink.clk
		.reset       (rst_controller_001_reset_out_reset)                                     //                    reset_sink.reset
	);

	nios2_secure_memory_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	nios2_secure_memory_led_pio led_pio (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_external_connection_export)       // external_connection.export
	);

	nios2_secure_memory_onchip_mem onchip_mem (
		.clk         (clk_clk),                                    //   clk1.clk
		.address     (mm_interconnect_1_onchip_mem_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_onchip_mem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_onchip_mem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_onchip_mem_s1_write),      //       .write
		.readdata    (mm_interconnect_1_onchip_mem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_onchip_mem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_onchip_mem_s1_byteenable), //       .byteenable
		.reset       (rst_controller_001_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req),     //       .reset_req
		.address2    (mm_interconnect_0_onchip_mem_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_mem_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_mem_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_mem_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_mem_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_mem_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_mem_s2_byteenable), //       .byteenable
		.clk2        (clk_clk),                                    //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),         // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req),     //       .reset_req
		.freeze      (1'b0)                                        // (terminated)
	);

	nios2_secure_memory_sys_clk_timer sys_clk_timer (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_1_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                       //   irq.irq
	);

	nios2_secure_memory_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) cpu_custom_instruction_master_translator (
		.ci_slave_dataa            (cpu_custom_instruction_master_dataa),                              //       ci_slave.dataa
		.ci_slave_datab            (cpu_custom_instruction_master_datab),                              //               .datab
		.ci_slave_result           (cpu_custom_instruction_master_result),                             //               .result
		.ci_slave_n                (cpu_custom_instruction_master_n),                                  //               .n
		.ci_slave_readra           (cpu_custom_instruction_master_readra),                             //               .readra
		.ci_slave_readrb           (cpu_custom_instruction_master_readrb),                             //               .readrb
		.ci_slave_writerc          (cpu_custom_instruction_master_writerc),                            //               .writerc
		.ci_slave_a                (cpu_custom_instruction_master_a),                                  //               .a
		.ci_slave_b                (cpu_custom_instruction_master_b),                                  //               .b
		.ci_slave_c                (cpu_custom_instruction_master_c),                                  //               .c
		.ci_slave_ipending         (cpu_custom_instruction_master_ipending),                           //               .ipending
		.ci_slave_estatus          (cpu_custom_instruction_master_estatus),                            //               .estatus
		.comb_ci_master_dataa      (cpu_custom_instruction_master_translator_comb_ci_master_dataa),    // comb_ci_master.dataa
		.comb_ci_master_datab      (cpu_custom_instruction_master_translator_comb_ci_master_datab),    //               .datab
		.comb_ci_master_result     (cpu_custom_instruction_master_translator_comb_ci_master_result),   //               .result
		.comb_ci_master_n          (cpu_custom_instruction_master_translator_comb_ci_master_n),        //               .n
		.comb_ci_master_readra     (cpu_custom_instruction_master_translator_comb_ci_master_readra),   //               .readra
		.comb_ci_master_readrb     (cpu_custom_instruction_master_translator_comb_ci_master_readrb),   //               .readrb
		.comb_ci_master_writerc    (cpu_custom_instruction_master_translator_comb_ci_master_writerc),  //               .writerc
		.comb_ci_master_a          (cpu_custom_instruction_master_translator_comb_ci_master_a),        //               .a
		.comb_ci_master_b          (cpu_custom_instruction_master_translator_comb_ci_master_b),        //               .b
		.comb_ci_master_c          (cpu_custom_instruction_master_translator_comb_ci_master_c),        //               .c
		.comb_ci_master_ipending   (cpu_custom_instruction_master_translator_comb_ci_master_ipending), //               .ipending
		.comb_ci_master_estatus    (cpu_custom_instruction_master_translator_comb_ci_master_estatus),  //               .estatus
		.ci_slave_multi_clk        (1'b0),                                                             //    (terminated)
		.ci_slave_multi_reset      (1'b0),                                                             //    (terminated)
		.ci_slave_multi_clken      (1'b0),                                                             //    (terminated)
		.ci_slave_multi_reset_req  (1'b0),                                                             //    (terminated)
		.ci_slave_multi_start      (1'b0),                                                             //    (terminated)
		.ci_slave_multi_done       (),                                                                 //    (terminated)
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                             //    (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                             //    (terminated)
		.ci_slave_multi_result     (),                                                                 //    (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                      //    (terminated)
		.ci_slave_multi_readra     (1'b0),                                                             //    (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                             //    (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                             //    (terminated)
		.ci_slave_multi_a          (5'b00000),                                                         //    (terminated)
		.ci_slave_multi_b          (5'b00000),                                                         //    (terminated)
		.ci_slave_multi_c          (5'b00000),                                                         //    (terminated)
		.multi_ci_master_clk       (),                                                                 //    (terminated)
		.multi_ci_master_reset     (),                                                                 //    (terminated)
		.multi_ci_master_clken     (),                                                                 //    (terminated)
		.multi_ci_master_reset_req (),                                                                 //    (terminated)
		.multi_ci_master_start     (),                                                                 //    (terminated)
		.multi_ci_master_done      (1'b0),                                                             //    (terminated)
		.multi_ci_master_dataa     (),                                                                 //    (terminated)
		.multi_ci_master_datab     (),                                                                 //    (terminated)
		.multi_ci_master_result    (32'b00000000000000000000000000000000),                             //    (terminated)
		.multi_ci_master_n         (),                                                                 //    (terminated)
		.multi_ci_master_readra    (),                                                                 //    (terminated)
		.multi_ci_master_readrb    (),                                                                 //    (terminated)
		.multi_ci_master_writerc   (),                                                                 //    (terminated)
		.multi_ci_master_a         (),                                                                 //    (terminated)
		.multi_ci_master_b         (),                                                                 //    (terminated)
		.multi_ci_master_c         ()                                                                  //    (terminated)
	);

	nios2_secure_memory_cpu_custom_instruction_master_comb_xconnect cpu_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (cpu_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (cpu_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (cpu_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (cpu_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (cpu_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (cpu_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (cpu_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (cpu_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (cpu_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (cpu_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (cpu_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (cpu_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (cpu_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (cpu_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (cpu_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (cpu_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (cpu_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) cpu_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (cpu_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (cpu_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (cpu_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (cpu_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (cpu_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (cpu_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (cpu_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                      // (terminated)
		.ci_master_readrb    (),                                                                      // (terminated)
		.ci_master_writerc   (),                                                                      // (terminated)
		.ci_master_a         (),                                                                      // (terminated)
		.ci_master_b         (),                                                                      // (terminated)
		.ci_master_c         (),                                                                      // (terminated)
		.ci_master_ipending  (),                                                                      // (terminated)
		.ci_master_estatus   (),                                                                      // (terminated)
		.ci_master_clk       (),                                                                      // (terminated)
		.ci_master_clken     (),                                                                      // (terminated)
		.ci_master_reset_req (),                                                                      // (terminated)
		.ci_master_reset     (),                                                                      // (terminated)
		.ci_master_start     (),                                                                      // (terminated)
		.ci_master_done      (1'b0),                                                                  // (terminated)
		.ci_slave_clk        (1'b0),                                                                  // (terminated)
		.ci_slave_clken      (1'b0),                                                                  // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                  // (terminated)
		.ci_slave_reset      (1'b0),                                                                  // (terminated)
		.ci_slave_start      (1'b0),                                                                  // (terminated)
		.ci_slave_done       ()                                                                       // (terminated)
	);

	nios2_secure_memory_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                         (clk_clk),                                                  //                                                       clk_0_clk.clk
		.custom_secure_mem_instructions_reset_sink_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                       // custom_secure_mem_instructions_reset_sink_reset_bridge_in_reset.reset
		.custom_secure_mem_instructions_avalon_master_address                  (custom_secure_mem_instructions_avalon_master_address),     //                    custom_secure_mem_instructions_avalon_master.address
		.custom_secure_mem_instructions_avalon_master_waitrequest              (custom_secure_mem_instructions_avalon_master_waitrequest), //                                                                .waitrequest
		.custom_secure_mem_instructions_avalon_master_byteenable               (custom_secure_mem_instructions_avalon_master_byteenable),  //                                                                .byteenable
		.custom_secure_mem_instructions_avalon_master_chipselect               (custom_secure_mem_instructions_avalon_master_chipselect),  //                                                                .chipselect
		.custom_secure_mem_instructions_avalon_master_readdata                 (custom_secure_mem_instructions_avalon_master_readdata),    //                                                                .readdata
		.custom_secure_mem_instructions_avalon_master_write                    (custom_secure_mem_instructions_avalon_master_write),       //                                                                .write
		.custom_secure_mem_instructions_avalon_master_writedata                (custom_secure_mem_instructions_avalon_master_writedata),   //                                                                .writedata
		.onchip_mem_s2_address                                                 (mm_interconnect_0_onchip_mem_s2_address),                  //                                                   onchip_mem_s2.address
		.onchip_mem_s2_write                                                   (mm_interconnect_0_onchip_mem_s2_write),                    //                                                                .write
		.onchip_mem_s2_readdata                                                (mm_interconnect_0_onchip_mem_s2_readdata),                 //                                                                .readdata
		.onchip_mem_s2_writedata                                               (mm_interconnect_0_onchip_mem_s2_writedata),                //                                                                .writedata
		.onchip_mem_s2_byteenable                                              (mm_interconnect_0_onchip_mem_s2_byteenable),               //                                                                .byteenable
		.onchip_mem_s2_chipselect                                              (mm_interconnect_0_onchip_mem_s2_chipselect),               //                                                                .chipselect
		.onchip_mem_s2_clken                                                   (mm_interconnect_0_onchip_mem_s2_clken)                     //                                                                .clken
	);

	nios2_secure_memory_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                               (clk_clk),                                                   //                             clk_0_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                            //       cpu_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // jtag_uart_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                     (cpu_data_master_address),                                   //                       cpu_data_master.address
		.cpu_data_master_waitrequest                 (cpu_data_master_waitrequest),                               //                                      .waitrequest
		.cpu_data_master_byteenable                  (cpu_data_master_byteenable),                                //                                      .byteenable
		.cpu_data_master_read                        (cpu_data_master_read),                                      //                                      .read
		.cpu_data_master_readdata                    (cpu_data_master_readdata),                                  //                                      .readdata
		.cpu_data_master_write                       (cpu_data_master_write),                                     //                                      .write
		.cpu_data_master_writedata                   (cpu_data_master_writedata),                                 //                                      .writedata
		.cpu_data_master_debugaccess                 (cpu_data_master_debugaccess),                               //                                      .debugaccess
		.cpu_instruction_master_address              (cpu_instruction_master_address),                            //                cpu_instruction_master.address
		.cpu_instruction_master_waitrequest          (cpu_instruction_master_waitrequest),                        //                                      .waitrequest
		.cpu_instruction_master_read                 (cpu_instruction_master_read),                               //                                      .read
		.cpu_instruction_master_readdata             (cpu_instruction_master_readdata),                           //                                      .readdata
		.cpu_instruction_master_readdatavalid        (cpu_instruction_master_readdatavalid),                      //                                      .readdatavalid
		.cpu_debug_mem_slave_address                 (mm_interconnect_1_cpu_debug_mem_slave_address),             //                   cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                   (mm_interconnect_1_cpu_debug_mem_slave_write),               //                                      .write
		.cpu_debug_mem_slave_read                    (mm_interconnect_1_cpu_debug_mem_slave_read),                //                                      .read
		.cpu_debug_mem_slave_readdata                (mm_interconnect_1_cpu_debug_mem_slave_readdata),            //                                      .readdata
		.cpu_debug_mem_slave_writedata               (mm_interconnect_1_cpu_debug_mem_slave_writedata),           //                                      .writedata
		.cpu_debug_mem_slave_byteenable              (mm_interconnect_1_cpu_debug_mem_slave_byteenable),          //                                      .byteenable
		.cpu_debug_mem_slave_waitrequest             (mm_interconnect_1_cpu_debug_mem_slave_waitrequest),         //                                      .waitrequest
		.cpu_debug_mem_slave_debugaccess             (mm_interconnect_1_cpu_debug_mem_slave_debugaccess),         //                                      .debugaccess
		.jtag_uart_avalon_jtag_slave_address         (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //           jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write           (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                      .write
		.jtag_uart_avalon_jtag_slave_read            (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                      .read
		.jtag_uart_avalon_jtag_slave_readdata        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                      .readdata
		.jtag_uart_avalon_jtag_slave_writedata       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                      .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                      .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect      (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                      .chipselect
		.led_pio_s1_address                          (mm_interconnect_1_led_pio_s1_address),                      //                            led_pio_s1.address
		.led_pio_s1_write                            (mm_interconnect_1_led_pio_s1_write),                        //                                      .write
		.led_pio_s1_readdata                         (mm_interconnect_1_led_pio_s1_readdata),                     //                                      .readdata
		.led_pio_s1_writedata                        (mm_interconnect_1_led_pio_s1_writedata),                    //                                      .writedata
		.led_pio_s1_chipselect                       (mm_interconnect_1_led_pio_s1_chipselect),                   //                                      .chipselect
		.onchip_mem_s1_address                       (mm_interconnect_1_onchip_mem_s1_address),                   //                         onchip_mem_s1.address
		.onchip_mem_s1_write                         (mm_interconnect_1_onchip_mem_s1_write),                     //                                      .write
		.onchip_mem_s1_readdata                      (mm_interconnect_1_onchip_mem_s1_readdata),                  //                                      .readdata
		.onchip_mem_s1_writedata                     (mm_interconnect_1_onchip_mem_s1_writedata),                 //                                      .writedata
		.onchip_mem_s1_byteenable                    (mm_interconnect_1_onchip_mem_s1_byteenable),                //                                      .byteenable
		.onchip_mem_s1_chipselect                    (mm_interconnect_1_onchip_mem_s1_chipselect),                //                                      .chipselect
		.onchip_mem_s1_clken                         (mm_interconnect_1_onchip_mem_s1_clken),                     //                                      .clken
		.sys_clk_timer_s1_address                    (mm_interconnect_1_sys_clk_timer_s1_address),                //                      sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                      (mm_interconnect_1_sys_clk_timer_s1_write),                  //                                      .write
		.sys_clk_timer_s1_readdata                   (mm_interconnect_1_sys_clk_timer_s1_readdata),               //                                      .readdata
		.sys_clk_timer_s1_writedata                  (mm_interconnect_1_sys_clk_timer_s1_writedata),              //                                      .writedata
		.sys_clk_timer_s1_chipselect                 (mm_interconnect_1_sys_clk_timer_s1_chipselect),             //                                      .chipselect
		.sysid_control_slave_address                 (mm_interconnect_1_sysid_control_slave_address),             //                   sysid_control_slave.address
		.sysid_control_slave_readdata                (mm_interconnect_1_sysid_control_slave_readdata)             //                                      .readdata
	);

	nios2_secure_memory_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
